
// (2) ʱ�� + ������ֵ
// md_sequential_blocking.v

module md_sequential_blocking(
    input clk,
    input IN_A,
    input IN_B,
    input IN_D,
    output OUT_A0,
    output reg [1:0] OUT_E
);

// 1. Variable Declaration (��������)
reg [1:0] c = 0;  // �� Verilog �У�reg ��������������ʱ����ʼֵ���� reg [1:0] c = 0;����������Ҫ���ڷ��棻�� FPGA �ۺ�ʱ����ʼֵͨ�������ԣ������� always ����ͨ����λ�߼����ó�ʼֵ��ȷ�����ۺ��ԡ�

// 2. Main Code (������)
always @(posedge clk) begin
    c = IN_A + IN_B;  // ������ֵ����˳��ִ�У������ɼ�ǰ�����
    OUT_E = c + IN_D;
end

// 3. Output Assignment (�����ֵ)
assign OUT_A0 = IN_A;

endmodule

