`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/11/16 15:50:27
// Design Name: 
// Module Name: db
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module db(
   input  wire clk,      // ϵͳʱ��
    input  wire sw,   // ��������
    output wire db        // ����������
);

    // ״̬����
    localparam [2:0]
        IDLE      = 3'b000,  // ����״̬
        PRESS_S1  = 3'b001,  // ����ȷ��״̬1
        PRESS_S2  = 3'b010,  // ����ȷ��״̬2
        PRESS_S3  = 3'b011,  // ����ȷ��״̬3
        PRESSED   = 3'b100,  // �����ȶ�״̬
        RELEASE_S1= 3'b101,  // �ͷ�ȷ��״̬1
        RELEASE_S2= 3'b110,  // �ͷ�ȷ��״̬2
        RELEASE_S3= 3'b111;  // �ͷ�ȷ��״̬3

    // ������λ��20λ@100MHzʱ�� �� 10ms��
    localparam CNT_WIDTH = 20;
    
    // �ڲ��źŶ���
    reg [2:0]            state_r = IDLE;  // ��ǰ״̬���ϵ��ʼ��ΪIDLE
    reg [2:0]            next_state;      // ��һ״̬
    reg [CNT_WIDTH-1:0]  count_r = 0;     // ���������ϵ��ʼ��Ϊ0
    wire                 time_up;          // ��ʱ��ɱ�־
    reg                  db_r;         // ����Ĵ���

    // �������߼�
    localparam MAX_COUNT = 20'hFFFFF;  // 20λȫ1
    assign time_up = (count_r == MAX_COUNT);
    
    always @(posedge clk) begin
        if (state_r != next_state)
            count_r <= 0;
        else if (count_r != MAX_COUNT)  // ��ֹ���
            count_r <= count_r + 1;
    end

    // ״̬�Ĵ���
    always @(posedge clk) begin
        state_r <= next_state;
    end

    // ״̬ת��������߼�
    always @(*) begin
        // Ĭ�ϱ��ֵ�ǰ״̬
        next_state = state_r;
        db_r = 1'b0;

        case (state_r)
            IDLE: begin
                if (sw)
                    next_state = PRESS_S1;
            end

            PRESS_S1: begin
                if (!sw)
                    next_state = IDLE;
                else if (time_up)
                    next_state = PRESS_S2;
            end

            PRESS_S2: begin
                if (!sw)
                    next_state = IDLE;
                else if (time_up)
                    next_state = PRESS_S3;
            end

            PRESS_S3: begin
                if (!sw)
                    next_state = IDLE;
                else if (time_up)
                    next_state = PRESSED;
            end

            PRESSED: begin
                db_r = 1'b1;
                if (!sw)
                    next_state = RELEASE_S1;
            end

            RELEASE_S1: begin
                db_r = 1'b1;
                if (sw)
                    next_state = PRESSED;
                else if (time_up)
                    next_state = RELEASE_S2;
            end

            RELEASE_S2: begin
                db_r = 1'b1;
                if (sw)
                    next_state = PRESSED;
                else if (time_up)
                    next_state = RELEASE_S3;
            end

            RELEASE_S3: begin
                db_r = 1'b1;
                if (sw)
                    next_state = PRESSED;
                else if (time_up)
                    next_state = IDLE;
            end

            default: next_state = IDLE;
        endcase
    end

    // �����ֵ
    assign db = db_r;

endmodule
